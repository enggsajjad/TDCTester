library verilog;
use verilog.vl_types.all;
entity tf2 is
end tf2;
