library verilog;
use verilog.vl_types.all;
entity tf is
end tf;
